module top_module( output one );

// Insert your code here
    assign one = 0;

endmodule
